module single_cycle_RISC-V(input clk ,rst);
	
endmodule
